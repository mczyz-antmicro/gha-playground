
module hello(input clk);

initial

begin: proc_he
	$display("helllo");
end

endmodule
